library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity vga_font is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic
);
end entity;

architecture prom of vga_font is
	type rom is array(0 to  16383) of std_logic;
	signal rom_data: rom := (
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','1','1','0','1','0','0','0','0','0','0','0','1','0',
		'1','0','0','0','0','0','0','0','1','0','0','0','0','0','1','0',
		'0','0','0','0','0','0','1','0','1','0','0','0','0','0','0','0',
		'1','0','0','0','0','0','1','0','0','0','0','0','0','0','1','0',
		'1','0','0','0','0','0','0','0','1','0','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','1','1','1','1','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','1','0','0','1','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','1','1','0','0','1','1','1','1','1','1','1','0',
		'0','1','1','0','1','1','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','1','1','0','0','1','1','1','1','1','1','1','0',
		'0','1','1','0','1','1','0','0','0','1','1','0','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','0','1','0','1','1','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','1','0','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','0','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','0','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','1','1','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','1','0','1','1','0','1','1','0','1','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','1','1','1','1','1','1','1','1',
		'0','0','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','1','1','1','1','1','1','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','0','0','1','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','1','0','0',
		'0','0','1','1','1','1','0','0','0','1','1','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','1','1','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','1','1','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','1','1','1','1','0','1','1','0','1','1','1','1','0',
		'1','1','0','1','1','1','1','0','1','1','0','1','1','1','0','0',
		'1','1','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','0','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'1','1','0','0','0','0','1','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','1','0',
		'0','1','1','0','0','1','1','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','1','1','1','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','0','1','0','0','1','1','0','1','0','0','0',
		'0','1','1','1','1','0','0','0','0','1','1','0','1','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','0','1','0','0','1','1','0','1','0','0','0',
		'0','1','1','1','1','0','0','0','0','1','1','0','1','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'1','1','0','0','0','0','1','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','1','1','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','0','1','1','1','0','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','1','1','1','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','1','1','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','1','1','0','0',
		'0','1','1','1','1','0','0','0','0','1','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','0','1','1','1','0',
		'1','1','1','1','1','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'1','1','1','1','0','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','0','1','1','1','1','0','1','1','0','0','1','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','1','1','1','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','1','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','1','1','1','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','1','1','1','0','0','1','1','1','1','1','1','0',
		'0','1','0','1','1','0','1','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','0','1','1','0','0',
		'0','0','1','1','1','0','0','0','0','0','0','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','1','0','1','1','1','0','0','1','1','0','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','0','1','1','1','1','1','0','0',
		'0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','1','1','1','0','0','0','1','1','0','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','1','1','1','1','0','1','1','0','0','0','1','1','0',
		'1','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','0','0','0','0','1','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','0','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','1','0','0','0','0','0',
		'0','1','1','1','0','0','0','0','0','0','1','1','1','0','0','0',
		'0','0','0','1','1','1','0','0','0','0','0','0','1','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','0','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','0','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','1',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','0','0','0',
		'0','0','0','0','1','1','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','1','1','1','1','0','0',
		'0','1','1','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'1','1','0','0','0','0','0','0','1','1','0','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','0','1','0','0','0','1','1','0','0','0','0','0',
		'1','1','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','0','1','1','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'0','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','1','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','1','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','1','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'1','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','0','1','1','1','1','0','0','0',
		'0','1','1','1','1','0','0','0','0','1','1','0','1','1','0','0',
		'0','1','1','0','0','1','1','0','1','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','1','0','1','1','0','0',
		'1','1','1','1','1','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','1','1','1','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','1','1','1','0','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','0','1','1','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','1','1','0','0','0','0','0','0','1','1','0','0',
		'0','0','0','1','1','1','1','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','1','1','1','0','0',
		'0','1','1','1','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','0','0','0','0','1','1','0','0','0','0','0',
		'0','1','1','0','0','0','0','0','1','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','1','1','1','0','0',
		'1','1','0','0','0','1','1','0','0','1','1','0','0','0','0','0',
		'0','0','1','1','1','0','0','0','0','0','0','0','1','1','0','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','1','1','1','1','1','1','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','0','0','0','0','0','1','1','0','0','0','0',
		'0','0','1','1','0','1','1','0','0','0','0','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','1','1','0','0','1','1','0','0',
		'1','1','0','0','1','1','0','0','0','1','1','1','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','1','1','0','0','1','1','0','0','1','1','0','0','1','1','0',
		'0','0','1','1','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','0','1','0','1','1','0','1','1','0','1','0','1','1','0',
		'1','1','1','1','1','1','1','0','0','1','1','0','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0',
		'0','1','1','0','1','1','0','0','0','0','1','1','1','0','0','0',
		'0','0','1','1','1','0','0','0','0','0','1','1','1','0','0','0',
		'0','1','1','0','1','1','0','0','1','1','0','0','0','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','1','1','0','0','0','1','1','0',
		'1','1','0','0','0','1','1','0','0','1','1','1','1','1','1','0',
		'0','0','0','0','0','1','1','0','0','0','0','0','1','1','0','0',
		'1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','1','1','1','1','1','1','1','0',
		'1','1','0','0','1','1','0','0','0','0','0','1','1','0','0','0',
		'0','0','1','1','0','0','0','0','0','1','1','0','0','0','0','0',
		'1','1','0','0','0','1','1','0','1','1','1','1','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','0','1','1','1','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','0','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','0','1','1','1','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','0','0','1','1','0','0','0',
		'0','0','0','1','1','0','0','0','0','1','1','1','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','1','1','1','0','1','1','0','1','1','0','1','1','1','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0',
		'0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0');
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
